`include "decoders.v"

module phi2(a, z);
  input [1:0] a;
  output [15:0] z;
  wire [3:0] y;

  decoder2_4 d_inst(.a(a), .z(y));
  assign z[0] = 1'b0;
  assign z[15] = 1'b1;

  assign z[5] = ~a[0];
  assign z[10] = a[0];
  assign z[3] = ~a[1];
  assign z[12] = a[1];

  assign z[1] = y[0];
  assign z[14] = ~y[0];
  assign z[2] = y[1];
  assign z[13] = ~y[1];
  assign z[4] = y[2];
  assign z[11] = ~y[2];
  assign z[8] = y[3];
  assign z[7] = ~y[3];

  assign z[3] = y[0] | y[1];
  assign z[12] = ~z[3];
  assign z[5] = y[0] | y[2];
  assign z[10] = ~z[5];
  assign z[9] = y[0] | y[3];
  assign z[6] = ~z[9];
  assign z[6] = y[1] | y[2];
  assign z[9] = ~z[6];
  assign z[10] = y[1] | y[3];
  assign z[5] = ~z[10];
  assign z[12] = y[2] | y[3];
  assign z[3] = ~z[12];
endmodule

module phi3(a, z);
  input [2:0] a;
  output [255:0] z;
  wire [7:0] y;

  decoder3_8 d_inst(.a(a), .z(y));
  assign z[0] = 1'b0;
  assign z[255] = 1'b1;

  assign z[85] = ~a[0];
  assign z[170] = a[0];
  assign z[51] = ~a[1];
  assign z[204] = a[1];
  assign z[15] = ~a[2];
  assign z[240] = a[2];

  assign z[1] = y[0];
  assign z[254] = ~y[0];
  assign z[2] = y[1];
  assign z[253] = ~y[1];
  assign z[4] = y[2];
  assign z[251] = ~y[2];
  assign z[8] = y[3];
  assign z[247] = ~y[3];
  assign z[16] = y[4];
  assign z[239] = ~y[4];
  assign z[32] = y[5];
  assign z[223] = ~y[5];
  assign z[64] = y[6];
  assign z[191] = ~y[6];
  assign z[128] = y[7];
  assign z[127] = ~y[7];

  assign z[3] = y[0] | y[1];
  assign z[252] = ~z[3];
  assign z[5] = y[0] | y[2];
  assign z[250] = ~z[5];
  assign z[9] = y[0] | y[3];
  assign z[246] = ~z[9];
  assign z[17] = y[0] | y[4];
  assign z[238] = ~z[17];
  assign z[33] = y[0] | y[5];
  assign z[222] = ~z[33];
  assign z[65] = y[0] | y[6];
  assign z[190] = ~z[65];
  assign z[129] = y[0] | y[7];
  assign z[126] = ~z[129];
  assign z[6] = y[1] | y[2];
  assign z[249] = ~z[6];
  assign z[10] = y[1] | y[3];
  assign z[245] = ~z[10];
  assign z[18] = y[1] | y[4];
  assign z[237] = ~z[18];
  assign z[34] = y[1] | y[5];
  assign z[221] = ~z[34];
  assign z[66] = y[1] | y[6];
  assign z[189] = ~z[66];
  assign z[130] = y[1] | y[7];
  assign z[125] = ~z[130];
  assign z[12] = y[2] | y[3];
  assign z[243] = ~z[12];
  assign z[20] = y[2] | y[4];
  assign z[235] = ~z[20];
  assign z[36] = y[2] | y[5];
  assign z[219] = ~z[36];
  assign z[68] = y[2] | y[6];
  assign z[187] = ~z[68];
  assign z[132] = y[2] | y[7];
  assign z[123] = ~z[132];
  assign z[24] = y[3] | y[4];
  assign z[231] = ~z[24];
  assign z[40] = y[3] | y[5];
  assign z[215] = ~z[40];
  assign z[72] = y[3] | y[6];
  assign z[183] = ~z[72];
  assign z[136] = y[3] | y[7];
  assign z[119] = ~z[136];
  assign z[48] = y[4] | y[5];
  assign z[207] = ~z[48];
  assign z[80] = y[4] | y[6];
  assign z[175] = ~z[80];
  assign z[144] = y[4] | y[7];
  assign z[111] = ~z[144];
  assign z[96] = y[5] | y[6];
  assign z[159] = ~z[96];
  assign z[160] = y[5] | y[7];
  assign z[95] = ~z[160];
  assign z[192] = y[6] | y[7];
  assign z[63] = ~z[192];

  assign z[7] = y[0] | z[6];
  assign z[248] = ~z[7];
  assign z[11] = y[0] | z[10];
  assign z[244] = ~z[11];
  assign z[19] = y[0] | z[18];
  assign z[236] = ~z[19];
  assign z[35] = y[0] | z[34];
  assign z[220] = ~z[35];
  assign z[67] = y[0] | z[66];
  assign z[188] = ~z[67];
  assign z[131] = y[0] | z[130];
  assign z[124] = ~z[131];
  assign z[13] = y[0] | z[12];
  assign z[242] = ~z[13];
  assign z[21] = y[0] | z[20];
  assign z[234] = ~z[21];
  assign z[37] = y[0] | z[36];
  assign z[218] = ~z[37];
  assign z[69] = y[0] | z[68];
  assign z[186] = ~z[69];
  assign z[133] = y[0] | z[132];
  assign z[122] = ~z[133];
  assign z[25] = y[0] | z[24];
  assign z[230] = ~z[25];
  assign z[41] = y[0] | z[40];
  assign z[214] = ~z[41];
  assign z[73] = y[0] | z[72];
  assign z[182] = ~z[73];
  assign z[137] = y[0] | z[136];
  assign z[118] = ~z[137];
  assign z[49] = y[0] | z[48];
  assign z[206] = ~z[49];
  assign z[81] = y[0] | z[80];
  assign z[174] = ~z[81];
  assign z[145] = y[0] | z[144];
  assign z[110] = ~z[145];
  assign z[97] = y[0] | z[96];
  assign z[158] = ~z[97];
  assign z[161] = y[0] | z[160];
  assign z[94] = ~z[161];
  assign z[193] = y[0] | z[192];
  assign z[62] = ~z[193];
  assign z[14] = y[1] | z[12];
  assign z[241] = ~z[14];
  assign z[22] = y[1] | z[20];
  assign z[233] = ~z[22];
  assign z[38] = y[1] | z[36];
  assign z[217] = ~z[38];
  assign z[70] = y[1] | z[68];
  assign z[185] = ~z[70];
  assign z[134] = y[1] | z[132];
  assign z[121] = ~z[134];
  assign z[26] = y[1] | z[24];
  assign z[229] = ~z[26];
  assign z[42] = y[1] | z[40];
  assign z[213] = ~z[42];
  assign z[74] = y[1] | z[72];
  assign z[181] = ~z[74];
  assign z[138] = y[1] | z[136];
  assign z[117] = ~z[138];
  assign z[50] = y[1] | z[48];
  assign z[205] = ~z[50];
  assign z[82] = y[1] | z[80];
  assign z[173] = ~z[82];
  assign z[146] = y[1] | z[144];
  assign z[109] = ~z[146];
  assign z[98] = y[1] | z[96];
  assign z[157] = ~z[98];
  assign z[162] = y[1] | z[160];
  assign z[93] = ~z[162];
  assign z[194] = y[1] | z[192];
  assign z[61] = ~z[194];
  assign z[28] = y[2] | z[24];
  assign z[227] = ~z[28];
  assign z[44] = y[2] | z[40];
  assign z[211] = ~z[44];
  assign z[76] = y[2] | z[72];
  assign z[179] = ~z[76];
  assign z[140] = y[2] | z[136];
  assign z[115] = ~z[140];
  assign z[52] = y[2] | z[48];
  assign z[203] = ~z[52];
  assign z[84] = y[2] | z[80];
  assign z[171] = ~z[84];
  assign z[148] = y[2] | z[144];
  assign z[107] = ~z[148];
  assign z[100] = y[2] | z[96];
  assign z[155] = ~z[100];
  assign z[164] = y[2] | z[160];
  assign z[91] = ~z[164];
  assign z[196] = y[2] | z[192];
  assign z[59] = ~z[196];
  assign z[56] = y[3] | z[48];
  assign z[199] = ~z[56];
  assign z[88] = y[3] | z[80];
  assign z[167] = ~z[88];
  assign z[152] = y[3] | z[144];
  assign z[103] = ~z[152];
  assign z[104] = y[3] | z[96];
  assign z[151] = ~z[104];
  assign z[168] = y[3] | z[160];
  assign z[87] = ~z[168];
  assign z[200] = y[3] | z[192];
  assign z[55] = ~z[200];
  assign z[112] = y[4] | z[96];
  assign z[143] = ~z[112];
  assign z[176] = y[4] | z[160];
  assign z[79] = ~z[176];
  assign z[208] = y[4] | z[192];
  assign z[47] = ~z[208];
  assign z[224] = y[5] | z[192];
  assign z[31] = ~z[224];

  assign z[23] = z[3] | z[20];
  assign z[232] = ~z[23];
  assign z[39] = z[3] | z[36];
  assign z[216] = ~z[39];
  assign z[71] = z[3] | z[68];
  assign z[184] = ~z[71];
  assign z[27] = z[3] | z[24];
  assign z[228] = ~z[27];
  assign z[43] = z[3] | z[40];
  assign z[212] = ~z[43];
  assign z[75] = z[3] | z[72];
  assign z[180] = ~z[75];
  assign z[83] = z[3] | z[80];
  assign z[172] = ~z[83];
  assign z[99] = z[3] | z[96];
  assign z[156] = ~z[99];
  assign z[29] = z[5] | z[24];
  assign z[226] = ~z[29];
  assign z[45] = z[5] | z[40];
  assign z[210] = ~z[45];
  assign z[77] = z[5] | z[72];
  assign z[178] = ~z[77];
  assign z[53] = z[5] | z[48];
  assign z[202] = ~z[53];
  assign z[101] = z[5] | z[96];
  assign z[154] = ~z[101];
  assign z[57] = z[9] | z[48];
  assign z[198] = ~z[57];
  assign z[89] = z[9] | z[80];
  assign z[166] = ~z[89];
  assign z[105] = z[9] | z[96];
  assign z[150] = ~z[105];
  assign z[113] = z[17] | z[96];
  assign z[142] = ~z[113];
  assign z[30] = z[6] | z[24];
  assign z[225] = ~z[30];
  assign z[46] = z[6] | z[40];
  assign z[209] = ~z[46];
  assign z[78] = z[6] | z[72];
  assign z[177] = ~z[78];
  assign z[54] = z[6] | z[48];
  assign z[201] = ~z[54];
  assign z[86] = z[6] | z[80];
  assign z[169] = ~z[86];
  assign z[102] = z[6] | z[96];
  assign z[153] = ~z[102];
  assign z[58] = z[10] | z[48];
  assign z[197] = ~z[58];
  assign z[90] = z[10] | z[80];
  assign z[165] = ~z[90];
  assign z[106] = z[10] | z[96];
  assign z[149] = ~z[106];
  assign z[114] = z[18] | z[96];
  assign z[141] = ~z[114];
  assign z[60] = z[12] | z[48];
  assign z[195] = ~z[60];
  assign z[92] = z[12] | z[80];
  assign z[163] = ~z[92];
  assign z[108] = z[12] | z[96];
  assign z[147] = ~z[108];
  assign z[116] = z[20] | z[96];
  assign z[139] = ~z[116];
  assign z[120] = z[24] | z[96];
  assign z[135] = ~z[120];
endmodule

